`ifndef MUL_MODEL_PKG
`define MUL_MODEL_PKG
package mul_model_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import mul_agent_pkg::*;
	`include "mul_model.sv"
endpackage
`endif
