`ifndef MUL_SEQ_LIST
`define MUL_SEQ_LIST
package mul_seq_list;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import mul_agent_pkg::*;
	import mul_model_pkg::*;
	import mul_env_pkg::*;

	`include "mul_basic_seq.sv"
endpackage
`endif
