`ifndef MUL_TEST_LIST
`define MUL_TEST_LIST
package mul_test_list;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	import mul_env_pkg::*;
	import mul_seq_list::*;

	`include "mul_basic_test.sv"

endpackage
`endif
