`define DWIDTH 8
`define NUM_TRANS 10
